library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

-- uMem interface
entity uMem is
  port (
    uAddr : in unsigned(12 downto 0);
    uData : out unsigned(31 downto 0));
end uMem;

architecture Behavioral of uMem is

-- micro Memory
type u_mem_t is array (0 to 42) of unsigned(31 downto 0);
constant u_mem_c : u_mem_t :=
   -- ALU_TB_FB_S_P_LC_SEQ_myADR
  (
   -- Hämtfas 00
   b"000_0011_0100_0_0_00_0000_0000000000000", -- ASR:=PC
   b"000_0010_0001_0_1_00_0000_0000000000000", -- IR:=PM, PC:=PC+1
   b"000_0000_0000_0_0_00_0010_0000000000000", -- uPC := K2
   
   -- Direktadressering 03
   b"000_0001_0100_0_0_00_0001_0000000000000", -- ASR:=IR, uPC:= K1
   
   -- Immediate 04
   b"000_0011_0100_0_1_00_0001_0000000000000", -- ASR:=PC, PC:= PC+1, uPC:= K1
   
   -- Indirekt adressering 05
   b"000_0001_0100_0_0_00_0000_0000000000000", -- ASR:= IR
   b"000_0010_0100_0_0_00_0001_0000000000000", -- ASR:= PM, uPC:= K1
   
   --Indexerad adressering 07
   b"001_0001_0000_0_0_00_0000_0000000000000", -- AR:= IR
   b"010_0110_0000_1_0_00_0000_0000000000000", -- AR:= GRX+AR
   b"000_0111_0100_1_0_00_0001_0000000000000", -- ASR:= AR, uPC:= K1
   
   -- Load 0A
   b"000_0010_0110_0_0_00_0011_0000000000000", -- Grx := PM(A)
   
   -- Store 0B
   b"000_0110_0010_0_0_00_0011_0000000000000", -- PM(A) := GRx
   
   -- Addi 0C
   b"001_0110_0000_0_0_00_0000_0000000000000", -- AR := GRx
   b"010_0010_0000_0_0_00_0000_0000000000000", -- AR := AR + PM(A)
   b"000_0111_0110_0_0_00_0011_0000000000000", -- GRx := AR
   
   -- SUBI 0F
   b"001_0110_0000_0_0_00_0000_0000000000000", -- AR := GRx
   b"011_0010_0000_0_0_00_0000_0000000000000", -- AR:= AR-PM
   b"000_0111_0110_0_0_00_0011_0000000000000", -- GRx := AR
   
   -- Andi 12
   b"001_0110_0000_0_0_00_0000_0000000000000", -- AR := GRx
   b"100_0010_0000_0_0_00_0000_0000000000000", -- AR := AR and PM(A)
   b"000_0111_0110_0_0_00_0011_0000000000000", -- GRx := AR
   
   -- GET_JOYSTICK 15
   b"000_1111_0110_0_0_00_0011_0000000000000", -- GRx := JOYSTICK
   
   -- Bra 16

   b"001_0011_0000_0_0_00_0000_0000000000000", -- AR := PC
   b"010_1000_0000_0_0_00_0000_0000000000000", -- AR += IR
   b"000_0111_0011_0_0_00_0011_0000000000000", -- PC := AR

  -- Bne 19
   b"000_0000_0000_0_0_00_0100_0000000010110", -- Om Z=0, hop xxxxxxx
   b"000_0000_0000_0_0_00_0011_0000000000000", -- Z=1
   
   -- Halt 1B
   b"000_0000_0000_0_0_00_1111_0000000000000", -- SEQ = 1111
   
   -- Cmpi 1C
   b"001_0010_0000_0_0_00_0000_0000000000000", -- AR := PM(A) 
   b"011_0110_0000_0_0_00_0011_0000000000000", -- AR -= GRx
   
   -- Bmi 1E
   b"000_0000_0000_0_0_00_1001_0000000010110", -- Om N=1 hopp BRA xxxxxxxx
   b"000_0000_0000_0_0_00_0011_0000000000000", -- else 00
   
   -- BGE 20
   b"000_0000_0000_0_0_00_1001_0000000100100", -- N=1, JMP 24 xxxxxx
   b"000_0000_0000_0_0_00_1011_0000000100100", -- V = 1, JMP 24
   b"000_0000_0000_0_0_00_0101_0000000010110", -- JMP BRA
   b"000_0000_0000_0_0_00_1011_0000000010110", -- V =1 JMP BRA
   b"000_0000_0000_0_0_00_0011_0000000000000", -- FINISH
  
   -- GET_RANDOM 25
   b"000_1001_0110_0_0_00_0011_0000000000000", -- Grx := out_reg_sync

   -- Beq 26
   b"000_0000_0000_0_0_00_1000_0000000010110", -- OM Z = 1, HOP xxxx
   b"000_0000_0000_0_0_00_0011_0000000000000",
   
   -- Ori 28
   b"001_0110_0000_0_0_00_0000_0000000000000", -- Ar := Grx
   b"101_0010_0000_0_0_00_0000_0000000000000", -- AR := AR | Pm(A)
   b"000_0111_0110_0_0_00_0011_0000000000000" -- Grx := AR
   );


begin  -- Behavioral
  uData <= u_mem_c(to_integer(uAddr));

end Behavioral;
